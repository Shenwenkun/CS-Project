`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2024/06/01 15:46:37
// Design Name: 
// Module Name: Bin2Hex
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Bin2Hex(
input clk,
input [3:0] bin_i,
output reg [7:0] segctrl_o
    );
    always @(posedge clk) begin
        case(bin_i)
        4'b0001:segctrl_o <= 8'b00001100;
        4'b0010:segctrl_o <= 8'b11011010;
        4'b0011:segctrl_o <= 8'b11110010;
        4'b0100:segctrl_o <= 8'b01100110;
        4'b0101:segctrl_o <= 8'b10110110;
        4'b0110:segctrl_o <= 8'b10111110;
        4'b0111:segctrl_o <= 8'b11100000;
        4'b1000:segctrl_o <= 8'b11111110;
        4'b1001:segctrl_o <= 8'b11110110;
        4'b1010:segctrl_o <= 8'b11101110;
        4'b1011:segctrl_o <= 8'b00111110;
        4'b1100:segctrl_o <= 8'b00011010;
        4'b1101:segctrl_o <= 8'b01111010;
        4'b1110:segctrl_o <= 8'b10011110;
        4'b1111:segctrl_o <= 8'b10001110;
        endcase
    end
endmodule
